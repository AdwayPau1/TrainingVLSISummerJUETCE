module half_subtractor(input a, b, output S, Cout);
//add your code here
endmodule
