module half_subtractor(input a, b, output reg S, Cout);
//your code here
endmodule
