module half_subtractor(input a, b, output D, B);
//your code here
endmodule
